`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Abhishek kumar
// 
// Create Date: 03.02.2025 20:26:09
// Design Name: 
// Module Name: two_one_mux
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module two_one_mux(
input [3:0]a,b,
input sel,
output reg [3:0]out
    );

always@(*)begin
    if(sel) out=b;
    else out=a;
end    
endmodule
